Pupusa de Maiz
nico
0 1 0
5 1 1 2 2 2 0 
3
0 0 4 67 5 150 
1 0 0 0 0 0 0 0 1 1 1 1 1 1 
0 7 9
